$dumpfile("dump.vcd");
$dumpvars;