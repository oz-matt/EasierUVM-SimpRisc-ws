`include "sequences/insgen_prand_ins_seq.sv"
`include "sequences/insgen_prand_inorder_ins_seq.sv"
