typedef enum {false, true} boolean;
