extern function init_params(boolean init_rx, instr_category_bm icbm);