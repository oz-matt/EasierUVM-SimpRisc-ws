import "DPI-C" function void get_reference_output(insgen_pkt_t ip);
export "DPI-C" function cpu_resolve;