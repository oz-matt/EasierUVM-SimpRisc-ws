instr_category_bm ibm = instr_category_bm'(STORE);

m_insgen_config.init_params(false, ibm);