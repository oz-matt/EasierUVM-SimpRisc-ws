
`include "tests/test_direct_ins.sv"
`include "tests/test_rand_ins.sv"
