import "DPI-C" function int something(insgen_pkt_t s);