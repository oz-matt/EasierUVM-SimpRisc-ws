
initial in_data_bus = 0;

/*clocking cb @(posedge clk);
	default input #2 output #2
	
endclocking*/