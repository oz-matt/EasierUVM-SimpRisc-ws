extern function void build_phase (uvm_phase phase);

uvm_blocking_get_port#(instruction_base_si) pull_port;
