
	extern function new(boolean init_rx, instr_category_bm icbm);
