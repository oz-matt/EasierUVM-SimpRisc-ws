instr_category_bm ibm = instr_category_bm'(LOAD | STORE | ARITHMETIC);

m_insgen_config.init_params(true, ibm);