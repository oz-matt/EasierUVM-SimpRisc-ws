typedef enum {false, true} boean;
