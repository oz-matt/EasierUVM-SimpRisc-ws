import "DPI-C" function void somethin(insgen_pkt_t ip);
export "DPI-C" function cpu_resolve;