extern task run_phase(uvm_phase phase);