
initial in_data_bus = 0;