$fsdbDumpfile("novas.fsdb");
$fsdbDumpvars();
$fsdbDumpon;
//$dumpfile("dump.vcd");
//$dumpvars;