constraint ins_c {
  instruction inside {32'h0040A003, 32'h00110113};
};
