import "DPI-C" function int something(int d);