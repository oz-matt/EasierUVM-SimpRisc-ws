
`include "tests/test_direct_ins.sv"
`include "tests/test_fill_cpu_rxs.sv"
