// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: _sequencer.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Fri Jul 10 01:43:41 2020
//=============================================================================
// Description: Sequencer for 
//=============================================================================

`ifndef _SEQUENCER_SV
`define _SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #() _sequencer_t;


`endif // _SEQUENCER_SV

