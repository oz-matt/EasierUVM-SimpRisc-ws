// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: memw_sequencer.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Tue Aug 18 07:39:50 2020
//=============================================================================
// Description: Sequencer for memw
//=============================================================================

`ifndef MEMW_SEQUENCER_SV
`define MEMW_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(memw_obj) memw_sequencer_t;


`endif // MEMW_SEQUENCER_SV

