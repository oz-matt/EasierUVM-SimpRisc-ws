
class rand_ins_gen extends uvm_component;
	
	//uvm_seq_item_pull_imp
	
	function new(string name, uvm_component parent);
		super.new(name, parent);
	endfunction
	
endclass
