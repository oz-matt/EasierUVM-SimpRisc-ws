
	typedef struct {
		arithmetic_instruction_si l;
		arithmetic_instruction_si a;
	} li_instruction_t;
	