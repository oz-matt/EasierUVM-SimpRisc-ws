function void reference::write_reference_0(trans_rand_ins t);
	`uvm_warning("P", $sformatf("In Ref!!: %s", t.ibsi.get_asm_string()))
endfunction