

// Each unique test must extend top_test and use a type override for a 
// sequence extended from insgen_default_seq
