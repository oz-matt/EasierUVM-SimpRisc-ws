// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: memr_sequencer.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Fri Jul 24 23:06:54 2020
//=============================================================================
// Description: Sequencer for memr
//=============================================================================

`ifndef MEMR_SEQUENCER_SV
`define MEMR_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(memr_obj) memr_sequencer_t;


`endif // MEMR_SEQUENCER_SV

