
	typedef struct {
		arithmetic_instruction_si l;
		arithmetic_instruction_si a;
	} li_instruction_t;
	
	
typedef struct {
	int instruction;
	int name;
} insgen_pkt_t;
