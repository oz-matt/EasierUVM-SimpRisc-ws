//tconfig = new;
