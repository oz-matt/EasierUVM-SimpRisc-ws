
class insgen_test_config;
	
	int init_cpu_regs_with_rand_vals;
	
	function new();
		init_cpu_regs_with_rand_vals = 1;
	endfunction
	
endclass
