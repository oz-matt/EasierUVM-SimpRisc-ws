insgen_test_config tconfig;

tconfig = new(true);
