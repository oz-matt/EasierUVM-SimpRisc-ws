rand_ins_gen rig;
