insgen_test_config tconfig;