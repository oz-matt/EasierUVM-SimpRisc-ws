// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: _if.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Fri Jul 10 01:43:41 2020
//=============================================================================
// Description: Signal interface for agent 
//=============================================================================

`ifndef _IF_SV
`define _IF_SV

interface (); 

  timeunit      1ns;
  timeprecision 1ps;

  import _pkg::*;


  // You can insert properties and assertions here

  // You can insert code here by setting if_inc_inside_interface in file 

endinterface : 

`endif // _IF_SV

