instruction_base_si isi[$];