// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: _pkg.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2017-01-19 on Fri Jul 10 01:43:41 2020
//=============================================================================
// Description: Package for agent 
//=============================================================================

package _pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;


  `include "_.sv"
  `include "_config.sv"
  `include "_driver.sv"
  `include "_monitor.sv"
  `include "_sequencer.sv"
  `include "_coverage.sv"
  `include "_agent.sv"
  `include "_seq_lib.sv"

endpackage : _pkg
