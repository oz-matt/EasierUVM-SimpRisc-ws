extern function void build_phase (uvm_phase phase);