uvm_seq_item_pull_port#(instruction_base_si) pull_port;
