extern function void start_of_simulation_phase(uvm_phase phase);