
package seq_ins_pkg;
	
	
	
endpackage
