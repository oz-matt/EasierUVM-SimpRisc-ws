//insgen_test_config tco;